module MAU
#(parameter matrix_dim = 8)
(
    input [7:0] host_instruction, data_in,
    input clk, reset,
    output wire  [7:0] data_out,
    output wire busy
);



endmodule