module Multiplier
#(parameter num_bits = 512)
(input  [num_bits-1:0] dd, aa,
input clk, reset,
output [num_bits-1:0] product,
output reg done_flag);

endmodule