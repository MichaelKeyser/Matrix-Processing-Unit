module Adder(input inbus1 , input i, input const, input const_flag, input start_flag, output reg done_flag);

endmodule