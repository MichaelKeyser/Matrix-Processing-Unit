module MAU
#(parameter matrix_dim = 8)
(
    input [7:0] host_instruction, data_in,
    input clk, reset,
    output [7:0] data_out,
    output busy_flag
);

endmodule